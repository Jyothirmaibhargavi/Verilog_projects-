module bcd_sevensegment_conv(D,a,b,c,d,e,f,g );
input[3:0]D;
output reg a,b,c,d,e,f,g;
 always @(*) 
 begin
 case(D)
 4'b0000: {a,b,c,d,e,f,g} = 7'b1111110;
 4'b0001: {a,b,c,d,e,f,g} = 7'b0110000;
 4'b0010: {a,b,c,d,e,f,g} = 7'b1101101;
 4'b0011: {a,b,c,d,e,f,g} = 7'b1111001;
 4'b0100: {a,b,c,d,e,f,g} = 7'b0110011;
 4'b0101: {a,b,c,d,e,f,g} = 7'b1011011;
 4'b0110: {a,b,c,d,e,f,g} = 7'b1011111;
 4'b0111: {a,b,c,d,e,f,g} = 7'b1110000;
 4'b1000: {a,b,c,d,e,f,g} = 7'b1111111;
 4'b1001: {a,b,c,d,e,f,g} = 7'b1111011;
 default: {a,b,c,d,e,f,g} = 7'b0000000;
 endcase
 end
endmodule

// Loading work.bcd_sevensegment_conv
//# a=1 b=1 c=1 d=1 e=1 f=1 g=0 D= 0
//# a=1 b=1 c=1 d=1 e=1 f=1 g=1 D= 8
//# a=1 b=1 c=1 d=0 e=0 f=0 g=0 D= 7
//# a=1 b=1 c=1 d=1 e=0 f=1 g=1 D= 9
//# a=0 b=0 c=0 d=0 e=0 f=0 g=0 D=12
